`ifndef sa_engine_ip_v1_0_tb_include_vh_
`define sa_engine_ip_v1_0_tb_include_vh_

//Configuration current bd names
`define BD_NAME sa_engine_ip_v1_0_bfm_1
`define BD_INST_NAME sa_engine_ip_v1_0_bfm_1_i
`define BD_WRAPPER sa_engine_ip_v1_0_bfm_1_wrapper

//Configuration address parameters

`endif

